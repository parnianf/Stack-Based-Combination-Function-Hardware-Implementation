library verilog;
use verilog.vl_types.all;
entity Comb_TB is
end Comb_TB;
